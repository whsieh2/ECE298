module brickMaker(input frame_clk, Reset,
					input logic[3:0] level,
					output logic[9:0] bX1, bY1, bX2, bY2, bX3, bY3, bX4, bY4, bX5, bY5, bX6, bY6, bX7, bY7, bX8, bY8, bX9, bY9, bX10, bY10, 
					bX11, bY11, bX12, bY12, bX13, bY13, bX14, bY14, bX15, bY15, bX16, bY16, bX17, bY17, bX18, bY18, bX19, bY19, bX20, bY20, 
					bX21, bY21, bX22, bY22, bX23, bY23, bX24, bY24, bX25, bY25, bX26, bY26, bX27, bY27, bX28, bY28, bX29, bY29, bX30, bY30, 
					bX31, bY31, bX32, bY32, bX33, bY33, bX34, bY34, bX35, bY35, bX36, bY36, bX37, bY37, bX38, bY38, bX39, bY39, bX40, bY40, 
					bX41, bY41, bX42, bY42, bX43, bY43, bX44, bY44, bX45, bY45, bX46, bY46, bX47, bY47, bX48, bY48, bX49, bY49, bX50, bY50, 
					bX51, bY51, bX52, bY52, bX53, bY53, bX54, bY54, bX55, bY55, bX56, bY56, bX57, bY57, bX58, bY58, bX59, bY59, bX60, bY60,
					bX61, bY61, bX62, bY62, bX63, bY63, bX64, bY64, bX65, bY65, bX66, bY66, bX67, bY67, bX68, bY68, bX69, bY69, bX70, bY70,
					bX71, bY71, bX72, bY72, bX73, bY73, bX74, bY74, bX75, bY75, bX76, bY76, bX77, bY77, bX78, bY78, bX79, bY79, bX80, bY80, 
					bX81, bY81, bX82, bY82, bX83, bY83, bX84, bY84, bX85, bY85, bX86, bY86, bX87, bY87, bX88, bY88, bX89, bY89, bX90, bY90, 
					bX91, bY91, bX92, bY92, bX93, bY93, bX94, bY94, bX95, bY95, bX96, bY96, bX97, bY97, bX98, bY98, bX99, bY99, bX100, bY100, 
					bX101, bY101, bX102, bY102, bX103, bY103, bX104, bY104, bX105, bY105, bX106, bY106, bX107, bY107, bX108, bY108, bX109, bY109, bX110, bY110,
					input logic [2:0]brick1, brick2, brick3, brick4,brick5,brick6,brick7,brick8,brick9,brick10,brick11,brick12,brick13,brick14,brick15,brick16,brick17,brick18,brick19,brick20,
					brick21, brick22, brick23, brick24,brick25,brick26,brick27,brick28,brick29,brick30,brick31,brick32,brick33,brick34,brick35,brick36,brick37,brick38,brick39,brick40,
					brick41, brick42, brick43, brick44,brick45,brick46,brick47,brick48,brick49,brick50,brick51,brick52,brick53,brick54,brick55,brick56,brick57,brick58,brick59,brick60,
					brick61, brick62, brick63, brick64,brick65,brick66,brick67,brick68,brick69,brick70,brick71,brick72,brick73,brick74,brick75,brick76,brick77,brick78,brick79,brick80,
					brick81,brick82,brick83,brick84,brick85,brick86,brick87,brick88,brick89,brick90,brick91,brick92,brick93,brick94,brick95,brick96,brick97,brick98,brick99,brick100,
					brick101,brick102,brick103,brick104,brick105,brick106,brick107,brick108,brick109,brick110,
					output logic[2:0] brickLevel_1, brickLevel_2, brickLevel_3, brickLevel_4,brickLevel_5,brickLevel_6,brickLevel_7,brickLevel_8,brickLevel_9,brickLevel_10,brickLevel_11,brickLevel_12,brickLevel_13,brickLevel_14,brickLevel_15,brickLevel_16,brickLevel_17,brickLevel_18,brickLevel_19,brickLevel_20,
					brickLevel_21, brickLevel_22, brickLevel_23, brickLevel_24,brickLevel_25,brickLevel_26,brickLevel_27,brickLevel_28,brickLevel_29,brickLevel_30,brickLevel_31,brickLevel_32,brickLevel_33,brickLevel_34,brickLevel_35,brickLevel_36,brickLevel_37,brickLevel_38,brickLevel_39,brickLevel_40,
					brickLevel_41, brickLevel_42, brickLevel_43, brickLevel_44,brickLevel_45,brickLevel_46,brickLevel_47,brickLevel_48,brickLevel_49,brickLevel_50,brickLevel_51,brickLevel_52,brickLevel_53,brickLevel_54,brickLevel_55,brickLevel_56,brickLevel_57,brickLevel_58,brickLevel_59,brickLevel_60,
					brickLevel_61, brickLevel_62, brickLevel_63, brickLevel_64,brickLevel_65,brickLevel_66,brickLevel_67,brickLevel_68,brickLevel_69,brickLevel_70,brickLevel_71, brickLevel_72, brickLevel_73, brickLevel_74,brickLevel_75,brickLevel_76,brickLevel_77,brickLevel_78,brickLevel_79,brickLevel_80,
					brickLevel_81,brickLevel_82,brickLevel_83,brickLevel_84,brickLevel_85,brickLevel_86,brickLevel_87,brickLevel_88,brickLevel_89,brickLevel_90,brickLevel_91, brickLevel_92, brickLevel_93, brickLevel_94,brickLevel_95,brickLevel_96,brickLevel_97,brickLevel_98,brickLevel_99,brickLevel_100,
					brickLevel_101,brickLevel_102,brickLevel_103,brickLevel_104,brickLevel_105,brickLevel_106,brickLevel_107,brickLevel_108,brickLevel_109,brickLevel_110);
// 0 > 217 Y each brick
// 0> 638 X each brick 57 
//Purple-> 3 lives (3'b111) -> 7 pts
//Yellow-> 2 lives (3'b101) -> 5 pts
//Orange-> 1 live  (3'b010) -> 2 pts
//Finishing a level -> 1 pt
always_ff //@ (posedge Reset or posedge frame_clk)
begin
	if (Reset)
	begin
		//Level 1, Score Before: 0, BrickScore:32,
		brickLevel_1<=3'b000;
		brickLevel_2<=3'b000;
		brickLevel_3<=3'b000;
		brickLevel_4<=3'b000;
		brickLevel_5<=3'b000;
		brickLevel_6<=3'b000;
		brickLevel_7<=3'b000;
		brickLevel_8<=3'b000;
		brickLevel_9<=3'b000;
		brickLevel_10<=3'b000;
		brickLevel_11<=3'b000;
		brickLevel_12<=3'b000;
		brickLevel_13<=3'b000;
		brickLevel_14<=3'b000;
		brickLevel_15<=3'b000;
		brickLevel_16<=3'b000;
		brickLevel_17<=3'b000;
		brickLevel_18<=3'b000;
		brickLevel_19<=3'b000;
		brickLevel_20<=3'b000;
		brickLevel_21<=3'b000;
		brickLevel_22<=3'b000;
		brickLevel_23<=3'b000;
		brickLevel_24<=3'b010;
		brickLevel_25<=3'b010;
		brickLevel_26<=3'b010;
		brickLevel_27<=3'b010;
		brickLevel_28<=3'b000;
		brickLevel_29<=3'b000;
		brickLevel_30<=3'b000;
		brickLevel_31<=3'b000;
		brickLevel_32<=3'b000;
		brickLevel_33<=3'b000;
		brickLevel_34<=3'b010;
		brickLevel_35<=3'b010;
		brickLevel_36<=3'b010;
		brickLevel_37<=3'b010;
		brickLevel_38<=3'b000;
		brickLevel_39<=3'b000;
		brickLevel_40<=3'b000;
		brickLevel_41<=3'b000;
		brickLevel_42<=3'b000;
		brickLevel_43<=3'b000;
		brickLevel_44<=3'b010;
		brickLevel_45<=3'b010;
		brickLevel_46<=3'b010;
		brickLevel_47<=3'b010;
		brickLevel_48<=3'b000;
		brickLevel_49<=3'b000;
		brickLevel_50<=3'b000;
		brickLevel_51<=3'b000;
		brickLevel_52<=3'b000;
		brickLevel_53<=3'b000;
		brickLevel_54<=3'b010;
		brickLevel_55<=3'b010;
		brickLevel_56<=3'b010;
		brickLevel_57<=3'b010;
		brickLevel_58<=3'b000;
		brickLevel_59<=3'b000;
		brickLevel_60<=3'b000;
		brickLevel_61<=3'b000;
		brickLevel_62<=3'b000;
		brickLevel_63<=3'b000;
		brickLevel_64<=3'b000;
		brickLevel_65<=3'b000;
		brickLevel_66<=3'b000;
		brickLevel_67<=3'b000;
		brickLevel_68<=3'b000;
		brickLevel_69<=3'b000;
		brickLevel_70<=3'b000;// After this should be 1/b0; for level 1
		brickLevel_71<=3'b000; 
		brickLevel_72<=3'b000; 
		brickLevel_73<=3'b000; 
		brickLevel_74<=3'b000;
		brickLevel_75<=3'b000;
		brickLevel_76<=3'b000;
		brickLevel_77<=3'b000;
		brickLevel_78<=3'b000;
		brickLevel_79<=3'b000;
		brickLevel_80<=3'b000;
		brickLevel_81<=3'b000;
		brickLevel_82<=3'b000;
		brickLevel_83<=3'b000;
		brickLevel_84<=3'b000;
		brickLevel_85<=3'b000;
		brickLevel_86<=3'b000;
		brickLevel_87<=3'b000;
		brickLevel_88<=3'b000;
		brickLevel_89<=3'b000;
		brickLevel_90<=3'b000;
		brickLevel_91<=3'b000; 
		brickLevel_92<=3'b000; 
		brickLevel_93<=3'b000; 
		brickLevel_94<=3'b000;
		brickLevel_95<=3'b000;
		brickLevel_96<=3'b000;
		brickLevel_97<=3'b000;
		brickLevel_98<=3'b000;
		brickLevel_99<=3'b000;
		brickLevel_100<=3'b000;
		brickLevel_101<=3'b000;
		brickLevel_102<=3'b000;
		brickLevel_103<=3'b000;
		brickLevel_104<=3'b000;
		brickLevel_105<=3'b000;
		brickLevel_106<=3'b000;
		brickLevel_107<=3'b000;
		brickLevel_108<=3'b000;
		brickLevel_109<=3'b000;
		brickLevel_110<=3'b000;
	
	end
	else if (level==4'b0001)//Level 2, Initial Score: 33, BrickScore:96,
	begin
		brickLevel_1<=3'b010;
		brickLevel_2<=3'b010;
		brickLevel_3<=3'b010;
		brickLevel_4<=3'b010;
		brickLevel_5<=3'b010;
		brickLevel_6<=3'b010;
		brickLevel_7<=3'b010;
		brickLevel_8<=3'b010;
		brickLevel_9<=3'b010;
		brickLevel_10<=3'b010;
		brickLevel_11<=3'b010;
		brickLevel_12<=3'b000;
		brickLevel_13<=3'b000;
		brickLevel_14<=3'b000;
		brickLevel_15<=3'b000;
		brickLevel_16<=3'b000;
		brickLevel_17<=3'b000;
		brickLevel_18<=3'b000;
		brickLevel_19<=3'b000;
		brickLevel_20<=3'b010;
		brickLevel_21<=3'b010;
		brickLevel_22<=3'b000;
		brickLevel_23<=3'b010;
		brickLevel_24<=3'b010;
		brickLevel_25<=3'b010;
		brickLevel_26<=3'b010;
		brickLevel_27<=3'b010;
		brickLevel_28<=3'b010;
		brickLevel_29<=3'b000;
		brickLevel_30<=3'b010;
		brickLevel_31<=3'b010;
		brickLevel_32<=3'b000;
		brickLevel_33<=3'b010;
		brickLevel_34<=3'b010;
		brickLevel_35<=3'b010;
		brickLevel_36<=3'b010;
		brickLevel_37<=3'b010;
		brickLevel_38<=3'b010;
		brickLevel_39<=3'b000;
		brickLevel_40<=3'b010;
		brickLevel_41<=3'b010;
		brickLevel_42<=3'b000;
		brickLevel_43<=3'b010;
		brickLevel_44<=3'b010;
		brickLevel_45<=3'b010;
		brickLevel_46<=3'b010;
		brickLevel_47<=3'b010;
		brickLevel_48<=3'b010;
		brickLevel_49<=3'b000;
		brickLevel_50<=3'b010;
		brickLevel_51<=3'b010;
		brickLevel_52<=3'b000;
		brickLevel_53<=3'b000;
		brickLevel_54<=3'b000;
		brickLevel_55<=3'b000;
		brickLevel_56<=3'b000;
		brickLevel_57<=3'b000;
		brickLevel_58<=3'b000;
		brickLevel_59<=3'b000;
		brickLevel_60<=3'b010;
		brickLevel_61<=3'b010;
		brickLevel_62<=3'b010;
		brickLevel_63<=3'b010;
		brickLevel_64<=3'b010;
		brickLevel_65<=3'b010;
		brickLevel_66<=3'b010;
		brickLevel_67<=3'b010;
		brickLevel_68<=3'b010;
		brickLevel_69<=3'b010;
		brickLevel_70<=3'b010;// After this should be 1/b0; for level 1
		brickLevel_71<=3'b000; 
		brickLevel_72<=3'b000; 
		brickLevel_73<=3'b000; 
		brickLevel_74<=3'b000;
		brickLevel_75<=3'b000;
		brickLevel_76<=3'b000;
		brickLevel_77<=3'b000;
		brickLevel_78<=3'b000;
		brickLevel_79<=3'b000;
		brickLevel_80<=3'b000;
		brickLevel_81<=3'b000;
		brickLevel_82<=3'b000;
		brickLevel_83<=3'b000;
		brickLevel_84<=3'b000;
		brickLevel_85<=3'b000;
		brickLevel_86<=3'b000;
		brickLevel_87<=3'b000;
		brickLevel_88<=3'b000;
		brickLevel_89<=3'b000;
		brickLevel_90<=3'b000;
		brickLevel_91<=3'b000; 
		brickLevel_92<=3'b000; 
		brickLevel_93<=3'b000; 
		brickLevel_94<=3'b000;
		brickLevel_95<=3'b000;
		brickLevel_96<=3'b000;
		brickLevel_97<=3'b000;
		brickLevel_98<=3'b000;
		brickLevel_99<=3'b000;
		brickLevel_100<=3'b000;
		brickLevel_101<=3'b000;
		brickLevel_102<=3'b000;
		brickLevel_103<=3'b000;
		brickLevel_104<=3'b000;
		brickLevel_105<=3'b000;
		brickLevel_106<=3'b000;
		brickLevel_107<=3'b000;
		brickLevel_108<=3'b000;
		brickLevel_109<=3'b000;
		brickLevel_110<=3'b000;
		
	end

		
	
	else if (level==4'b0010)//Level 3, Initial Score: 97, BrickScore:96,
	begin
	brickLevel_1<=3'b111;
	brickLevel_2<=3'b000;
	brickLevel_3<=3'b000;
	brickLevel_4<=3'b000;
	brickLevel_5<=3'b111;
	brickLevel_6<=3'b000;
	brickLevel_7<=3'b000;
	brickLevel_8<=3'b000;
	brickLevel_9<=3'b111;
	brickLevel_10<=3'b000;
	brickLevel_11<=3'b000;
	brickLevel_12<=3'b101;
	brickLevel_13<=3'b000;
	brickLevel_14<=3'b101;
	brickLevel_15<=3'b000;
	brickLevel_16<=3'b101;
	brickLevel_17<=3'b000;
	brickLevel_18<=3'b101;
	brickLevel_19<=3'b000;
	brickLevel_20<=3'b101;
	brickLevel_21<=3'b000;
	brickLevel_22<=3'b000;
	brickLevel_23<=3'b010;
	brickLevel_24<=3'b000;
	brickLevel_25<=3'b000;
	brickLevel_26<=3'b000;
	brickLevel_27<=3'b010;
	brickLevel_28<=3'b000;
	brickLevel_29<=3'b000;
	brickLevel_30<=3'b000;
	brickLevel_31<=3'b000;
	brickLevel_32<=3'b101;
	brickLevel_33<=3'b000;
	brickLevel_34<=3'b101;
	brickLevel_35<=3'b000;
	brickLevel_36<=3'b101;
	brickLevel_37<=3'b000;
	brickLevel_38<=3'b101;
	brickLevel_39<=3'b000;
	brickLevel_40<=3'b101;
	brickLevel_41<=3'b111;
	brickLevel_42<=3'b000;
	brickLevel_43<=3'b000;
	brickLevel_44<=3'b000;
	brickLevel_45<=3'b111;
	brickLevel_46<=3'b000;
	brickLevel_47<=3'b000;
	brickLevel_48<=3'b000;
	brickLevel_49<=3'b111;
	brickLevel_50<=3'b000;
	brickLevel_51<=3'b000;
	brickLevel_52<=3'b000;
	brickLevel_53<=3'b000;
	brickLevel_54<=3'b000;
	brickLevel_55<=3'b000;
	brickLevel_56<=3'b000;
	brickLevel_57<=3'b000;
	brickLevel_58<=3'b000;
	brickLevel_59<=3'b000;
	brickLevel_60<=3'b000;
	brickLevel_61<=3'b000;
	brickLevel_62<=3'b000;
	brickLevel_63<=3'b000;
	brickLevel_64<=3'b000;
	brickLevel_65<=3'b000;
	brickLevel_66<=3'b000;
	brickLevel_67<=3'b000;
	brickLevel_68<=3'b000;
	brickLevel_69<=3'b000;
	brickLevel_70<=3'b000;// After this should be 1/b0; for level 1
	brickLevel_71<=3'b000; 
	brickLevel_72<=3'b000; 
	brickLevel_73<=3'b000; 
	brickLevel_74<=3'b000;
	brickLevel_75<=3'b000;
	brickLevel_76<=3'b000;
	brickLevel_77<=3'b000;
	brickLevel_78<=3'b000;
	brickLevel_79<=3'b000;
	brickLevel_80<=3'b000;
	brickLevel_81<=3'b000;
	brickLevel_82<=3'b000;
	brickLevel_83<=3'b000;
	brickLevel_84<=3'b000;
	brickLevel_85<=3'b000;
	brickLevel_86<=3'b000;
	brickLevel_87<=3'b000;
	brickLevel_88<=3'b000;
	brickLevel_89<=3'b000;
	brickLevel_90<=3'b000;
	brickLevel_91<=3'b000; 
	brickLevel_92<=3'b000; 
	brickLevel_93<=3'b000; 
	brickLevel_94<=3'b000;
	brickLevel_95<=3'b000;
	brickLevel_96<=3'b000;
	brickLevel_97<=3'b000;
	brickLevel_98<=3'b000;
	brickLevel_99<=3'b000;
	brickLevel_100<=3'b000;
	brickLevel_101<=3'b000;
	brickLevel_102<=3'b000;
	brickLevel_103<=3'b000;
	brickLevel_104<=3'b000;
	brickLevel_105<=3'b000;
	brickLevel_106<=3'b000;
	brickLevel_107<=3'b000;
	brickLevel_108<=3'b000;
	brickLevel_109<=3'b000;
	brickLevel_110<=3'b000;
	
	end

else if (level==4'b0011)//Level 4, Initial Score: 194, BrickScore:247,
	begin
	//level<=4'b0011;
	brickLevel_1<=3'b111;
	brickLevel_2<=3'b111;
	brickLevel_3<=3'b111;
	brickLevel_4<=3'b101;
	brickLevel_5<=3'b101;
	brickLevel_6<=3'b101;
	brickLevel_7<=3'b101;
	brickLevel_8<=3'b111;
	brickLevel_9<=3'b111;
	brickLevel_10<=3'b111;
	brickLevel_11<=3'b111;
	brickLevel_12<=3'b000;
	brickLevel_13<=3'b000;
	brickLevel_14<=3'b101;
	brickLevel_15<=3'b000;
	brickLevel_16<=3'b000;
	brickLevel_17<=3'b000;
	brickLevel_18<=3'b111;
	brickLevel_19<=3'b000;
	brickLevel_20<=3'b000;
	brickLevel_21<=3'b111;
	brickLevel_22<=3'b000;
	brickLevel_23<=3'b000;
	brickLevel_24<=3'b101;
	brickLevel_25<=3'b000;
	brickLevel_26<=3'b000;
	brickLevel_27<=3'b000;
	brickLevel_28<=3'b111;
	brickLevel_29<=3'b000;
	brickLevel_30<=3'b000;
	brickLevel_31<=3'b111;
	brickLevel_32<=3'b111;
	brickLevel_33<=3'b111;
	brickLevel_34<=3'b101;
	brickLevel_35<=3'b000;
	brickLevel_36<=3'b000;
	brickLevel_37<=3'b000;
	brickLevel_38<=3'b111;
	brickLevel_39<=3'b111;
	brickLevel_40<=3'b111;
	brickLevel_41<=3'b111;
	brickLevel_42<=3'b000;
	brickLevel_43<=3'b000;
	brickLevel_44<=3'b101;
	brickLevel_45<=3'b000;
	brickLevel_46<=3'b000;
	brickLevel_47<=3'b000;
	brickLevel_48<=3'b111;
	brickLevel_49<=3'b000;
	brickLevel_50<=3'b000;
	brickLevel_51<=3'b111;
	brickLevel_52<=3'b000;
	brickLevel_53<=3'b000;
	brickLevel_54<=3'b101;
	brickLevel_55<=3'b000;
	brickLevel_56<=3'b000;
	brickLevel_57<=3'b000;
	brickLevel_58<=3'b111;
	brickLevel_59<=3'b000;
	brickLevel_60<=3'b000;
	brickLevel_61<=3'b111;
	brickLevel_62<=3'b111;
	brickLevel_63<=3'b111;
	brickLevel_64<=3'b101;
	brickLevel_65<=3'b101;
	brickLevel_66<=3'b101;
	brickLevel_67<=3'b101;
	brickLevel_68<=3'b111;
	brickLevel_69<=3'b111;
	brickLevel_70<=3'b111;// After this should be 1/b0; for level 1
	brickLevel_71<=3'b000; 
	brickLevel_72<=3'b000; 
	brickLevel_73<=3'b000; 
	brickLevel_74<=3'b000;
	brickLevel_75<=3'b000;
	brickLevel_76<=3'b000;
	brickLevel_77<=3'b000;
	brickLevel_78<=3'b000;
	brickLevel_79<=3'b000;
	brickLevel_80<=3'b000;
	brickLevel_81<=3'b000;
	brickLevel_82<=3'b000;
	brickLevel_83<=3'b000;
	brickLevel_84<=3'b000;
	brickLevel_85<=3'b000;
	brickLevel_86<=3'b000;
	brickLevel_87<=3'b000;
	brickLevel_88<=3'b000;
	brickLevel_89<=3'b000;
	brickLevel_90<=3'b000;
	brickLevel_91<=3'b000; 
	brickLevel_92<=3'b000; 
	brickLevel_93<=3'b000; 
	brickLevel_94<=3'b000;
	brickLevel_95<=3'b000;
	brickLevel_96<=3'b000;
	brickLevel_97<=3'b000;
	brickLevel_98<=3'b000;
	brickLevel_99<=3'b000;
	brickLevel_100<=3'b000;
	brickLevel_101<=3'b000;
	brickLevel_102<=3'b000;
	brickLevel_103<=3'b000;
	brickLevel_104<=3'b000;
	brickLevel_105<=3'b000;
	brickLevel_106<=3'b000;
	brickLevel_107<=3'b000;
	brickLevel_108<=3'b000;
	brickLevel_109<=3'b000;
	brickLevel_110<=3'b000;
	
	end
	else if (level==4'b0100)//Level 5, Initial Score: 442, BrickScore:194
	begin
	brickLevel_1<=3'b111;
	brickLevel_2<=3'b111;
	brickLevel_3<=3'b111;
	brickLevel_4<=3'b010;
	brickLevel_5<=3'b010;
	brickLevel_6<=3'b010;
	brickLevel_7<=3'b101;
	brickLevel_8<=3'b101;
	brickLevel_9<=3'b101;
	brickLevel_10<=3'b000;
	brickLevel_11<=3'b000;
	brickLevel_12<=3'b000;
	brickLevel_13<=3'b111;
	brickLevel_14<=3'b010;
	brickLevel_15<=3'b000;
	brickLevel_16<=3'b010;
	brickLevel_17<=3'b101;
	brickLevel_18<=3'b000;
	brickLevel_19<=3'b000;
	brickLevel_20<=3'b000;
	brickLevel_21<=3'b000;
	brickLevel_22<=3'b000;
	brickLevel_23<=3'b111;
	brickLevel_24<=3'b010;
	brickLevel_25<=3'b000;
	brickLevel_26<=3'b010;
	brickLevel_27<=3'b101;
	brickLevel_28<=3'b000;
	brickLevel_29<=3'b000;
	brickLevel_30<=3'b000;
	brickLevel_31<=3'b111;
	brickLevel_32<=3'b111;
	brickLevel_33<=3'b111;
	brickLevel_34<=3'b010;
	brickLevel_35<=3'b010;
	brickLevel_36<=3'b010;
	brickLevel_37<=3'b101;
	brickLevel_38<=3'b101;
	brickLevel_39<=3'b101;
	brickLevel_40<=3'b000;
	brickLevel_41<=3'b000;
	brickLevel_42<=3'b000;
	brickLevel_43<=3'b111;
	brickLevel_44<=3'b010;
	brickLevel_45<=3'b000;
	brickLevel_46<=3'b010;
	brickLevel_47<=3'b000;
	brickLevel_48<=3'b000;
	brickLevel_49<=3'b000;
	brickLevel_50<=3'b101;
	brickLevel_51<=3'b000;
	brickLevel_52<=3'b000;
	brickLevel_53<=3'b111;
	brickLevel_54<=3'b010;
	brickLevel_55<=3'b000;
	brickLevel_56<=3'b010;
	brickLevel_57<=3'b101;
	brickLevel_58<=3'b000;
	brickLevel_59<=3'b000;
	brickLevel_60<=3'b101;
	brickLevel_61<=3'b111;
	brickLevel_62<=3'b111;
	brickLevel_63<=3'b111;
	brickLevel_64<=3'b010;
	brickLevel_65<=3'b010;
	brickLevel_66<=3'b010;
	brickLevel_67<=3'b000;
	brickLevel_68<=3'b101;
	brickLevel_69<=3'b101;
	brickLevel_70<=3'b000;// After this should be 1/b0; for level 1
	brickLevel_71<=3'b000; 
	brickLevel_72<=3'b000; 
	brickLevel_73<=3'b000; 
	brickLevel_74<=3'b000;
	brickLevel_75<=3'b000;
	brickLevel_76<=3'b000;
	brickLevel_77<=3'b000;
	brickLevel_78<=3'b000;
	brickLevel_79<=3'b000;
	brickLevel_80<=3'b000;
	brickLevel_81<=3'b000;
	brickLevel_82<=3'b000;
	brickLevel_83<=3'b000;
	brickLevel_84<=3'b000;
	brickLevel_85<=3'b000;
	brickLevel_86<=3'b000;
	brickLevel_87<=3'b000;
	brickLevel_88<=3'b000;
	brickLevel_89<=3'b000;
	brickLevel_90<=3'b000;
	brickLevel_91<=3'b000; 
	brickLevel_92<=3'b000; 
	brickLevel_93<=3'b000; 
	brickLevel_94<=3'b000;
	brickLevel_95<=3'b000;
	brickLevel_96<=3'b000;
	brickLevel_97<=3'b000;
	brickLevel_98<=3'b000;
	brickLevel_99<=3'b000;
	brickLevel_100<=3'b000;
	brickLevel_101<=3'b000;
	brickLevel_102<=3'b000;
	brickLevel_103<=3'b000;
	brickLevel_104<=3'b000;
	brickLevel_105<=3'b000;
	brickLevel_106<=3'b000;
	brickLevel_107<=3'b000;
	brickLevel_108<=3'b000;
	brickLevel_109<=3'b000;
	brickLevel_110<=3'b000;
	
	end

else if (level==4'b0101)//Level 6, Initial Score: 637, BrickScore:134,
	begin
	brickLevel_1<=3'b111;
	brickLevel_2<=3'b111;
	brickLevel_3<=3'b111;
	brickLevel_4<=3'b111;
	brickLevel_5<=3'b111;
	brickLevel_6<=3'b111;
	brickLevel_7<=3'b111;
	brickLevel_8<=3'b111;
	brickLevel_9<=3'b111;
	brickLevel_10<=3'b111;
	brickLevel_11<=3'b000;
	brickLevel_12<=3'b101;
	brickLevel_13<=3'b101;
	brickLevel_14<=3'b101;
	brickLevel_15<=3'b101;
	brickLevel_16<=3'b101;
	brickLevel_17<=3'b101;
	brickLevel_18<=3'b101;
	brickLevel_19<=3'b101;
	brickLevel_20<=3'b000;
	brickLevel_21<=3'b000;
	brickLevel_22<=3'b000;
	brickLevel_23<=3'b010;
	brickLevel_24<=3'b010;
	brickLevel_25<=3'b010;
	brickLevel_26<=3'b010;
	brickLevel_27<=3'b010;
	brickLevel_28<=3'b010;
	brickLevel_29<=3'b000;
	brickLevel_30<=3'b000;
	brickLevel_31<=3'b000;
	brickLevel_32<=3'b000;
	brickLevel_33<=3'b000;
	brickLevel_34<=3'b010;
	brickLevel_35<=3'b010;
	brickLevel_36<=3'b010;
	brickLevel_37<=3'b010;
	brickLevel_38<=3'b000;
	brickLevel_39<=3'b000;
	brickLevel_40<=3'b000;
	brickLevel_41<=3'b000;
	brickLevel_42<=3'b000;
	brickLevel_43<=3'b000;
	brickLevel_44<=3'b000;
	brickLevel_45<=3'b010;
	brickLevel_46<=3'b010;
	brickLevel_47<=3'b000;
	brickLevel_48<=3'b000;
	brickLevel_49<=3'b000;
	brickLevel_50<=3'b000;
	brickLevel_51<=3'b000;
	brickLevel_52<=3'b000;
	brickLevel_53<=3'b000;
	brickLevel_54<=3'b000;
	brickLevel_55<=3'b000;
	brickLevel_56<=3'b000;
	brickLevel_57<=3'b000;
	brickLevel_58<=3'b000;
	brickLevel_59<=3'b000;
	brickLevel_60<=3'b000;
	brickLevel_61<=3'b000;
	brickLevel_62<=3'b000;
	brickLevel_63<=3'b000;
	brickLevel_64<=3'b000;
	brickLevel_65<=3'b000;
	brickLevel_66<=3'b000;
	brickLevel_67<=3'b000;
	brickLevel_68<=3'b000;
	brickLevel_69<=3'b000;
	brickLevel_70<=3'b000;
	brickLevel_71<=3'b000; 
	brickLevel_72<=3'b000; 
	brickLevel_73<=3'b000; 
	brickLevel_74<=3'b000;
	brickLevel_75<=3'b000;
	brickLevel_76<=3'b000;
	brickLevel_77<=3'b000;
	brickLevel_78<=3'b000;
	brickLevel_79<=3'b000;
	brickLevel_80<=3'b000;
	brickLevel_81<=3'b000;
	brickLevel_82<=3'b000;
	brickLevel_83<=3'b000;
	brickLevel_84<=3'b000;
	brickLevel_85<=3'b000;
	brickLevel_86<=3'b000;
	brickLevel_87<=3'b000;
	brickLevel_88<=3'b000;
	brickLevel_89<=3'b000;
	brickLevel_90<=3'b000;
	brickLevel_91<=3'b000; 
	brickLevel_92<=3'b000; 
	brickLevel_93<=3'b000; 
	brickLevel_94<=3'b000;
	brickLevel_95<=3'b000;
	brickLevel_96<=3'b000;
	brickLevel_97<=3'b000;
	brickLevel_98<=3'b000;
	brickLevel_99<=3'b000;
	brickLevel_100<=3'b000;
	brickLevel_101<=3'b000;
	brickLevel_102<=3'b000;
	brickLevel_103<=3'b000;
	brickLevel_104<=3'b000;
	brickLevel_105<=3'b000;
	brickLevel_106<=3'b000;
	brickLevel_107<=3'b000;
	brickLevel_108<=3'b000;
	brickLevel_109<=3'b000;
	brickLevel_110<=3'b000;

	end


else if (level==4'b0110)//Level 7, Initial Score: 772, BrickScore:246,
	begin
	brickLevel_1<=3'b000;
	brickLevel_2<=3'b111;
	brickLevel_3<=3'b010;
	brickLevel_4<=3'b010;
	brickLevel_5<=3'b010;
	brickLevel_6<=3'b010;
	brickLevel_7<=3'b010;
	brickLevel_8<=3'b010;
	brickLevel_9<=3'b111;
	brickLevel_10<=3'b000;
	brickLevel_11<=3'b101;
	brickLevel_12<=3'b000;
	brickLevel_13<=3'b111;
	brickLevel_14<=3'b010;
	brickLevel_15<=3'b010;
	brickLevel_16<=3'b010;
	brickLevel_17<=3'b010;
	brickLevel_18<=3'b111;
	brickLevel_19<=3'b000;
	brickLevel_20<=3'b101;
	brickLevel_21<=3'b010;
	brickLevel_22<=3'b101;
	brickLevel_23<=3'b000;
	brickLevel_24<=3'b111;
	brickLevel_25<=3'b010;
	brickLevel_26<=3'b010;
	brickLevel_27<=3'b111;
	brickLevel_28<=3'b000;
	brickLevel_29<=3'b101;
	brickLevel_30<=3'b010;
	brickLevel_31<=3'b010;
	brickLevel_32<=3'b010;
	brickLevel_33<=3'b101;
	brickLevel_34<=3'b000;
	brickLevel_35<=3'b111;
	brickLevel_36<=3'b111;
	brickLevel_37<=3'b000;
	brickLevel_38<=3'b101;
	brickLevel_39<=3'b010;
	brickLevel_40<=3'b010;
	brickLevel_41<=3'b101;
	brickLevel_42<=3'b101;
	brickLevel_43<=3'b101;
	brickLevel_44<=3'b101;
	brickLevel_45<=3'b000;
	brickLevel_46<=3'b000;
	brickLevel_47<=3'b101;
	brickLevel_48<=3'b101;
	brickLevel_49<=3'b101;
	brickLevel_50<=3'b101;
	brickLevel_51<=3'b000;
	brickLevel_52<=3'b000;
	brickLevel_53<=3'b000;
	brickLevel_54<=3'b000;
	brickLevel_55<=3'b111;
	brickLevel_56<=3'b111;
	brickLevel_57<=3'b000;
	brickLevel_58<=3'b000;
	brickLevel_59<=3'b000;
	brickLevel_60<=3'b000;
	brickLevel_61<=3'b000;
	brickLevel_62<=3'b000;
	brickLevel_63<=3'b000;
	brickLevel_64<=3'b000;
	brickLevel_65<=3'b000;
	brickLevel_66<=3'b000;
	brickLevel_67<=3'b000;
	brickLevel_68<=3'b000;
	brickLevel_69<=3'b000;
	brickLevel_70<=3'b000;// After this should be 1/b0; for level 1
	brickLevel_71<=3'b000; 
	brickLevel_72<=3'b000; 
	brickLevel_73<=3'b000; 
	brickLevel_74<=3'b000;
	brickLevel_75<=3'b000;
	brickLevel_76<=3'b000;
	brickLevel_77<=3'b000;
	brickLevel_78<=3'b000;
	brickLevel_79<=3'b000;
	brickLevel_80<=3'b000;
	brickLevel_81<=3'b000;
	brickLevel_82<=3'b000;
	brickLevel_83<=3'b000;
	brickLevel_84<=3'b000;
	brickLevel_85<=3'b000;
	brickLevel_86<=3'b000;
	brickLevel_87<=3'b000;
	brickLevel_88<=3'b000;
	brickLevel_89<=3'b000;
	brickLevel_90<=3'b000;
	brickLevel_91<=3'b000; 
	brickLevel_92<=3'b000; 
	brickLevel_93<=3'b000; 
	brickLevel_94<=3'b000;
	brickLevel_95<=3'b000;
	brickLevel_96<=3'b000;
	brickLevel_97<=3'b000;
	brickLevel_98<=3'b000;
	brickLevel_99<=3'b000;
	brickLevel_100<=3'b000;
	brickLevel_101<=3'b000;
	brickLevel_102<=3'b000;
	brickLevel_103<=3'b000;
	brickLevel_104<=3'b000;
	brickLevel_105<=3'b000;
	brickLevel_106<=3'b000;
	brickLevel_107<=3'b000;
	brickLevel_108<=3'b000;
	brickLevel_109<=3'b000;
	brickLevel_110<=3'b000;
	
	end

	else if (level==4'b0111)//Level 8, Initial Score: 1023, BrickScore:364, Total~: 1568
	begin
	brickLevel_1<=3'b111;
	brickLevel_2<=3'b111;
	brickLevel_3<=3'b111;
	brickLevel_4<=3'b101;
	brickLevel_5<=3'b101;
	brickLevel_6<=3'b101;
	brickLevel_7<=3'b101;
	brickLevel_8<=3'b111;
	brickLevel_9<=3'b111;
	brickLevel_10<=3'b111;
	brickLevel_11<=3'b101;
	brickLevel_12<=3'b101;
	brickLevel_13<=3'b101;
	brickLevel_14<=3'b010;
	brickLevel_15<=3'b010;
	brickLevel_16<=3'b010;
	brickLevel_17<=3'b010;
	brickLevel_18<=3'b101;
	brickLevel_19<=3'b101;
	brickLevel_20<=3'b101;
	brickLevel_21<=3'b111;
	brickLevel_22<=3'b000;
	brickLevel_23<=3'b000;
	brickLevel_24<=3'b010;
	brickLevel_25<=3'b010;
	brickLevel_26<=3'b010;
	brickLevel_27<=3'b010;
	brickLevel_28<=3'b000;
	brickLevel_29<=3'b000;
	brickLevel_30<=3'b000;
	brickLevel_31<=3'b000;
	brickLevel_32<=3'b000;
	brickLevel_33<=3'b000;
	brickLevel_34<=3'b010;
	brickLevel_35<=3'b010;
	brickLevel_36<=3'b010;
	brickLevel_37<=3'b010;
	brickLevel_38<=3'b000;
	brickLevel_39<=3'b000;
	brickLevel_40<=3'b111;
	brickLevel_41<=3'b111;
	brickLevel_42<=3'b111;
	brickLevel_43<=3'b111;
	brickLevel_44<=3'b111;
	brickLevel_45<=3'b111;
	brickLevel_46<=3'b111;
	brickLevel_47<=3'b111;
	brickLevel_48<=3'b111;
	brickLevel_49<=3'b111;
	brickLevel_50<=3'b111;
	brickLevel_51<=3'b000;
	brickLevel_52<=3'b010;
	brickLevel_53<=3'b000;
	brickLevel_54<=3'b010;
	brickLevel_55<=3'b000;
	brickLevel_56<=3'b000;
	brickLevel_57<=3'b010;
	brickLevel_58<=3'b000;
	brickLevel_59<=3'b010;
	brickLevel_60<=3'b000;
	brickLevel_61<=3'b010;
	brickLevel_62<=3'b000;
	brickLevel_63<=3'b010;
	brickLevel_64<=3'b000;
	brickLevel_65<=3'b010;
	brickLevel_66<=3'b010;
	brickLevel_67<=3'b000;
	brickLevel_68<=3'b010;
	brickLevel_69<=3'b000;
	brickLevel_70<=3'b010;
	brickLevel_71<=3'b111; 
	brickLevel_72<=3'b111; 
	brickLevel_73<=3'b111; 
	brickLevel_74<=3'b111;
	brickLevel_75<=3'b111;
	brickLevel_76<=3'b111;
	brickLevel_77<=3'b111;
	brickLevel_78<=3'b111;
	brickLevel_79<=3'b111;
	brickLevel_80<=3'b101;
	brickLevel_81<=3'b101;
	brickLevel_82<=3'b101;
	brickLevel_83<=3'b101;
	brickLevel_84<=3'b101;
	brickLevel_85<=3'b101;
	brickLevel_86<=3'b101;
	brickLevel_87<=3'b101;
	brickLevel_88<=3'b101;
	brickLevel_89<=3'b101;
	brickLevel_90<=3'b101;
	brickLevel_91<=3'b010; 
	brickLevel_92<=3'b010; 
	brickLevel_93<=3'b010; 
	brickLevel_94<=3'b010;
	brickLevel_95<=3'b010;
	brickLevel_96<=3'b010;
	brickLevel_97<=3'b010;
	brickLevel_98<=3'b010;
	brickLevel_99<=3'b010;
	brickLevel_100<=3'b000;
	brickLevel_101<=3'b000;
	brickLevel_102<=3'b000;
	brickLevel_103<=3'b000;
	brickLevel_104<=3'b000;
	brickLevel_105<=3'b000;
	brickLevel_106<=3'b000;
	brickLevel_107<=3'b000;
	brickLevel_108<=3'b000;
	brickLevel_109<=3'b000;
	brickLevel_110<=3'b000;
	
	end
	else//(level==4'b1000)//End Game Module
	begin
	brickLevel_1<=3'b111;
	brickLevel_2<=3'b111;
	brickLevel_3<=3'b111;
	brickLevel_4<=3'b101;
	brickLevel_5<=3'b000;
	brickLevel_6<=3'b000;
	brickLevel_7<=3'b101;
	brickLevel_8<=3'b010;
	brickLevel_9<=3'b010;
	brickLevel_10<=3'b000;
	
	brickLevel_11<=3'b111;
	brickLevel_12<=3'b000;
	brickLevel_13<=3'b000;
	brickLevel_14<=3'b101;
	brickLevel_15<=3'b101;
	brickLevel_16<=3'b000;
	brickLevel_17<=3'b101;
	brickLevel_18<=3'b010;
	brickLevel_19<=3'b000;
	brickLevel_20<=3'b010;
	
	brickLevel_21<=3'b111;
	brickLevel_22<=3'b111;
	brickLevel_23<=3'b111;
	brickLevel_24<=3'b101;
	brickLevel_25<=3'b000;
	brickLevel_26<=3'b101;
	brickLevel_27<=3'b101;
	brickLevel_28<=3'b010;
	brickLevel_29<=3'b000;
	brickLevel_30<=3'b010;
	
	brickLevel_31<=3'b111;
	brickLevel_32<=3'b000;
	brickLevel_33<=3'b000;
	brickLevel_34<=3'b101;
	brickLevel_35<=3'b000;
	brickLevel_36<=3'b000;
	brickLevel_37<=3'b101;
	brickLevel_38<=3'b010;
	brickLevel_39<=3'b000;
	brickLevel_40<=3'b010;
	
	brickLevel_41<=3'b111;
	brickLevel_42<=3'b111;
	brickLevel_43<=3'b111;
	brickLevel_44<=3'b101;
	brickLevel_45<=3'b000;
	brickLevel_46<=3'b000;
	brickLevel_47<=3'b101;
	brickLevel_48<=3'b010;
	brickLevel_49<=3'b010;
	brickLevel_50<=3'b000;
	
	brickLevel_51<=3'b000;
	brickLevel_52<=3'b000;
	brickLevel_53<=3'b000;
	brickLevel_54<=3'b000;
	brickLevel_55<=3'b000;
	brickLevel_56<=3'b000;
	brickLevel_57<=3'b000;
	brickLevel_58<=3'b000;
	brickLevel_59<=3'b000;
	brickLevel_60<=3'b000;
	
	brickLevel_61<=3'b000;
	brickLevel_62<=3'b000;
	brickLevel_63<=3'b000;
	brickLevel_64<=3'b000;
	brickLevel_65<=3'b000;
	brickLevel_66<=3'b000;
	brickLevel_67<=3'b000;
	brickLevel_68<=3'b000;
	brickLevel_69<=3'b000;
	brickLevel_70<=3'b000;// After this should be 1/b0; for level 1
	brickLevel_71<=3'b000; 
	brickLevel_72<=3'b000; 
	brickLevel_73<=3'b000; 
	brickLevel_74<=3'b000;
	brickLevel_75<=3'b000;
	brickLevel_76<=3'b000;
	brickLevel_77<=3'b000;
	brickLevel_78<=3'b000;
	brickLevel_79<=3'b000;
	brickLevel_80<=3'b000;
	brickLevel_81<=3'b000;
	brickLevel_82<=3'b000;
	brickLevel_83<=3'b000;
	brickLevel_84<=3'b000;
	brickLevel_85<=3'b000;
	brickLevel_86<=3'b000;
	brickLevel_87<=3'b000;
	brickLevel_88<=3'b000;
	brickLevel_89<=3'b000;
	brickLevel_90<=3'b000;
	brickLevel_91<=3'b000; 
	brickLevel_92<=3'b000; 
	brickLevel_93<=3'b000; 
	brickLevel_94<=3'b000;
	brickLevel_95<=3'b000;
	brickLevel_96<=3'b000;
	brickLevel_97<=3'b000;
	brickLevel_98<=3'b000;
	brickLevel_99<=3'b000;
	brickLevel_100<=3'b000;
	brickLevel_101<=3'b000;
	brickLevel_102<=3'b000;
	brickLevel_103<=3'b000;
	brickLevel_104<=3'b000;
	brickLevel_105<=3'b000;
	brickLevel_106<=3'b000;
	brickLevel_107<=3'b000;
	brickLevel_108<=3'b000;
	brickLevel_109<=3'b000;
	brickLevel_110<=3'b000;
	
	end
end
always_comb
begin
		bX1<=3;
		bY1<=4;
		bY2<=4;
		bX2<=66;
		bY3<=4;
		bX3<=129;
		bY4<=4;
		bX4<=192;
		bY5<=4;
		bX5<=255;
		bY6<=4;
		bX6<=318;
		bY7<=4;
		bX7<=381;
		bY8<=4;
		bX8<=444;
		bY9<=4;
		bX9<=507;
		bY10<=4;
		bX10<=570;
		
		bY11<=20;
		bX11<=3;
		bY12<=20;
		bX12<=66;
		bY13<=20;
		bX13<=129;
		bY14<=20;
		bX14<=192;
		bY15<=20;
		bX15<=255;
		bY16<=20;
		bX16<=318;
		bY17<=20;
		bX17<=381;
		bY18<=20;
		bX18<=444;
		bY19<=20;
		bX19<=507;
		bY20<=20;
		bX20<=570;
			
		bY21<=36;
		bX21<=3;
		bY22<=36;
		bX22<=66;
		bY23<=36;
		bX23<=129;
		bY24<=36;
		bX24<=192;
		bY25<=36;
		bX25<=255;
		bY26<=36;
		bX26<=318;
		bY27<=36;
		bX27<=381;
		bY28<=36;
		bX28<=444;
		bY29<=36;
		bX29<=507;
		bY30<=36;
		bX30<=570;
		
		bY31<=52;
		bX31<=3;
		bY32<=52;
		bX32<=66;
		bY33<=52;
		bX33<=129;
		bY34<=52;
		bX34<=192;
		bX35<=255;
		bY35<=52;
		bX36<=318;
		bY36<=52;
		bX37<=381;
		bY37<=52;
		bX38<=444;
		bY38<=52;
		bX39<=507;
		bY39<=52;
		bX40<=570;
		bY40<=52;
		
		bX41<=3;
		bY41<=68;
		bX42<=66;
		bY42<=68;
		bX43<=129;
		bY43<=68;
		bX44<=192;
		bY44<=68;
		bX45<=255;
		bY45<=68;
		bX46<=318;
		bY46<=68;
		bX47<=381;
		bY47<=68;
		bX48<=444;
		bY48<=68;
		bX49<=507;
		bY49<=68;
		bX50<=570;
		bY50<=68;
		
		bX51<=3;
		bY51<=84;
		bX52<=66;
		bY52<=84;
		bX53<=129;
		bY53<=84;
		bX54<=192;
		bY54<=84;
		bX55<=255;
		bY55<=84;
		bX56<=318;
		bY56<=84;
		bX57<=381;
		bY57<=84;
		bX58<=444;
		bY58<=84;
		bX59<=507;
		bY59<=84;
		bX60<=570;
		bY60<=84;
				
		bX61<=3;
		bY61<=100;
		bX62<=66;
		bY62<=100;
		bX63<=129;
		bY63<=100;
		bX64<=192;
		bY64<=100;
		bX65<=255;
		bY65<=100;
		bX66<=318;
		bY66<=100;
		bX67<=381;
		bY67<=100;
		bX68<=444;
		bY68<=100;
		bX69<=507;
		bY69<=100;
		bX70<=570;
		bY70<=100;
		
		bX71<=3;
		bY71<=116;
		bX72<=66;
		bY72<=116;
		bX73<=129;
		bY73<=116;
		bX74<=192;
		bY74<=116;
		bX75<=255;
		bY75<=116;
		bX76<=318;
		bY76<=116;
		bX77<=381;
		bY77<=116;
		bX78<=444;
		bY78<=116;
		bX79<=507;
		bY79<=116;
		bX80<=570;
		bY80<=116;
		
		bX81<=3;
		bY81<=132;
		bX82<=66;
		bY82<=132;
		bX83<=129;
		bY83<=132;
		bX84<=192;
		bY84<=132;
		bX85<=255;
		bY85<=132;
		bX86<=318;
		bY86<=132;
		bX87<=381;
		bY87<=132;
		bX88<=444;
		bY88<=132;
		bX89<=507;
		bY89<=132;
		bX90<=570;
		bY90<=132;
		
		bX91<=3;
		bY91<=148;
		bX92<=66;
		bY92<=148;
		bX93<=129;
		bY93<=148;
		bX94<=192;
		bY94<=148;
		bX95<=255;
		bY95<=148;
		bX96<=318;
		bY96<=148;
		bX97<=381;
		bY97<=148;
		bX98<=444;
		bY98<=148;
		bX99<=507;
		bY99<=148;
		bX100<=570;
		bY100<=148;
		
		bX101<=3;
		bY101<=164;
		bX102<=66;
		bY102<=164;
		bX103<=129;
		bY103<=164;
		bX104<=192;
		bY104<=164;
		bX105<=255;
		bY105<=164;
		bX106<=318;
		bY106<=164;
		bX107<=381;
		bY107<=164;
		bX108<=444;
		bY108<=164;
		bX109<=507;
		bY109<=164;
		bX110<=570;
		bY110<=164;
	end
endmodule
