module InvMixColumns_128 ( input[127:0] in,
						output logic [127:0] out );
					 
					 
InvMixColumns InMuxColumns0(.in(in[31:0]),.out(out[31:0]));
InvMixColumns InMuxColumns1(.in(in[63:32]),.out(out[63:32]));
InvMixColumns InMuxColumns2(.in(in[95:64]),.out(out[95:64]));
InvMixColumns InMuxColumns3(.in(in[127:96]),.out(out[127:96]));

endmodule